*ac sim command for cable impedance measurement
*lumped transmission line model with 20 segments per meter at 50 meters
*and a 50.000000 meter long cable
*one 10cm segment for a lumped transmission line model

*copyright � 2021 <analog devices>
*permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the �software�), to deal in the software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the software, and to permit persons to whom the software is furnished to do so, subject to the following conditions:
*the above copyright notice and this permission notice shall be included in all copies or substantial portions of the software.
*the software is provided �as is�, without warranty of any kind, express or implied, including but not limited to the warranties of merchantability, fitness for a particular purpose and noninfringement. in no event shall the authors or copyright holders be liable for any claim, damages or other liability, whether in an action of contract, tort or otherwise, arising from, out of or in connection with the software or the use or other dealings in the software.


.subckt tlump t1p t1n t2p t2n rtn
rx t1p rtn 1e9
g1 t1p a t1p a laplace=1/(1.134268e-5*((abs(s)/(2*pi))^0.5))
l1 a t2p {1*20.6435n}
c1 t2p rtn {1*2.25026p}
r1 t1n rtn 1e-6
r2 t2n rtn 1e-6
.ends tlump
*simple pd model for transmission line simulations

*copyright � 2021 <analog devices>
*permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the �software�), to deal in the software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the software, and to permit persons to whom the software is furnished to do so, subject to the following conditions:
*the above copyright notice and this permission notice shall be included in all copies or substantial portions of the software.
*the software is provided �as is�, without warranty of any kind, express or implied, including but not limited to the warranties of merchantability, fitness for a particular purpose and noninfringement. in no event shall the authors or copyright holders be liable for any claim, damages or other liability, whether in an action of contract, tort or otherwise, arising from, out of or in connection with the software or the use or other dealings in the software.


.subckt pd p n 0
*lpodl p n 80e-6
cpodl p n 15p
rpodl p n 10k
.ends pd
.param clump=1.6675e-12
.param llump=1.6675e-08
.param rg=100e6
.param rser=0.188
xseg0000 p0000 n0000 p0001 n0001 0 tlump
xseg0001 p0001 n0001 p0002 n0002 0 tlump
xseg0002 p0002 n0002 p0003 n0003 0 tlump
xseg0003 p0003 n0003 p0004 n0004 0 tlump
xseg0004 p0004 n0004 p0005 n0005 0 tlump
xseg0005 p0005 n0005 p0006 n0006 0 tlump
xseg0006 p0006 n0006 p0007 n0007 0 tlump
xseg0007 p0007 n0007 p0008 n0008 0 tlump
xseg0008 p0008 n0008 p0009 n0009 0 tlump
xseg0009 p0009 n0009 p0010 n0010 0 tlump
xseg0010 p0010 n0010 p0011 n0011 0 tlump
xseg0011 p0011 n0011 p0012 n0012 0 tlump
xseg0012 p0012 n0012 p0013 n0013 0 tlump
xseg0013 p0013 n0013 p0014 n0014 0 tlump
xseg0014 p0014 n0014 p0015 n0015 0 tlump
xseg0015 p0015 n0015 p0016 n0016 0 tlump
xseg0016 p0016 n0016 p0017 n0017 0 tlump
xseg0017 p0017 n0017 p0018 n0018 0 tlump
xseg0018 p0018 n0018 p0019 n0019 0 tlump
xseg0019 p0019 n0019 p0020 n0020 0 tlump
xseg0020 p0020 n0020 p0021 n0021 0 tlump
xseg0021 p0021 n0021 p0022 n0022 0 tlump
xseg0022 p0022 n0022 p0023 n0023 0 tlump
xseg0023 p0023 n0023 p0024 n0024 0 tlump
xseg0024 p0024 n0024 p0025 n0025 0 tlump
xseg0025 p0025 n0025 p0026 n0026 0 tlump
xseg0026 p0026 n0026 p0027 n0027 0 tlump
xseg0027 p0027 n0027 p0028 n0028 0 tlump
xseg0028 p0028 n0028 p0029 n0029 0 tlump
xseg0029 p0029 n0029 p0030 n0030 0 tlump
xseg0030 p0030 n0030 p0031 n0031 0 tlump
xseg0031 p0031 n0031 p0032 n0032 0 tlump
xseg0032 p0032 n0032 p0033 n0033 0 tlump
xseg0033 p0033 n0033 p0034 n0034 0 tlump
xseg0034 p0034 n0034 p0035 n0035 0 tlump
xseg0035 p0035 n0035 p0036 n0036 0 tlump
xseg0036 p0036 n0036 p0037 n0037 0 tlump
xseg0037 p0037 n0037 p0038 n0038 0 tlump
xseg0038 p0038 n0038 p0039 n0039 0 tlump
xseg0039 p0039 n0039 p0040 n0040 0 tlump
xseg0040 p0040 n0040 p0041 n0041 0 tlump
xseg0041 p0041 n0041 p0042 n0042 0 tlump
xseg0042 p0042 n0042 p0043 n0043 0 tlump
xseg0043 p0043 n0043 p0044 n0044 0 tlump
xseg0044 p0044 n0044 p0045 n0045 0 tlump
xseg0045 p0045 n0045 p0046 n0046 0 tlump
xseg0046 p0046 n0046 p0047 n0047 0 tlump
xseg0047 p0047 n0047 p0048 n0048 0 tlump
xseg0048 p0048 n0048 p0049 n0049 0 tlump
xseg0049 p0049 n0049 p0050 n0050 0 tlump
xseg0050 p0050 n0050 p0051 n0051 0 tlump
xseg0051 p0051 n0051 p0052 n0052 0 tlump
xseg0052 p0052 n0052 p0053 n0053 0 tlump
xseg0053 p0053 n0053 p0054 n0054 0 tlump
xseg0054 p0054 n0054 p0055 n0055 0 tlump
xseg0055 p0055 n0055 p0056 n0056 0 tlump
xseg0056 p0056 n0056 p0057 n0057 0 tlump
xseg0057 p0057 n0057 p0058 n0058 0 tlump
xseg0058 p0058 n0058 p0059 n0059 0 tlump
xseg0059 p0059 n0059 p0060 n0060 0 tlump
xseg0060 p0060 n0060 p0061 n0061 0 tlump
xseg0061 p0061 n0061 p0062 n0062 0 tlump
xseg0062 p0062 n0062 p0063 n0063 0 tlump
xseg0063 p0063 n0063 p0064 n0064 0 tlump
xseg0064 p0064 n0064 p0065 n0065 0 tlump
xseg0065 p0065 n0065 p0066 n0066 0 tlump
xseg0066 p0066 n0066 p0067 n0067 0 tlump
xseg0067 p0067 n0067 p0068 n0068 0 tlump
xseg0068 p0068 n0068 p0069 n0069 0 tlump
xseg0069 p0069 n0069 p0070 n0070 0 tlump
xseg0070 p0070 n0070 p0071 n0071 0 tlump
xseg0071 p0071 n0071 p0072 n0072 0 tlump
xseg0072 p0072 n0072 p0073 n0073 0 tlump
xseg0073 p0073 n0073 p0074 n0074 0 tlump
xseg0074 p0074 n0074 p0075 n0075 0 tlump
xseg0075 p0075 n0075 p0076 n0076 0 tlump
xseg0076 p0076 n0076 p0077 n0077 0 tlump
xseg0077 p0077 n0077 p0078 n0078 0 tlump
xseg0078 p0078 n0078 p0079 n0079 0 tlump
xseg0079 p0079 n0079 p0080 n0080 0 tlump
xseg0080 p0080 n0080 p0081 n0081 0 tlump
xseg0081 p0081 n0081 p0082 n0082 0 tlump
xseg0082 p0082 n0082 p0083 n0083 0 tlump
xseg0083 p0083 n0083 p0084 n0084 0 tlump
xseg0084 p0084 n0084 p0085 n0085 0 tlump
xseg0085 p0085 n0085 p0086 n0086 0 tlump
xseg0086 p0086 n0086 p0087 n0087 0 tlump
xseg0087 p0087 n0087 p0088 n0088 0 tlump
xseg0088 p0088 n0088 p0089 n0089 0 tlump
xseg0089 p0089 n0089 p0090 n0090 0 tlump
xseg0090 p0090 n0090 p0091 n0091 0 tlump
xseg0091 p0091 n0091 p0092 n0092 0 tlump
xseg0092 p0092 n0092 p0093 n0093 0 tlump
xseg0093 p0093 n0093 p0094 n0094 0 tlump
xseg0094 p0094 n0094 p0095 n0095 0 tlump
xseg0095 p0095 n0095 p0096 n0096 0 tlump
xseg0096 p0096 n0096 p0097 n0097 0 tlump
xseg0097 p0097 n0097 p0098 n0098 0 tlump
xseg0098 p0098 n0098 p0099 n0099 0 tlump
xseg0099 p0099 n0099 p0100 n0100 0 tlump
xseg0100 p0100 n0100 p0101 n0101 0 tlump
xseg0101 p0101 n0101 p0102 n0102 0 tlump
xseg0102 p0102 n0102 p0103 n0103 0 tlump
xseg0103 p0103 n0103 p0104 n0104 0 tlump
xseg0104 p0104 n0104 p0105 n0105 0 tlump
xseg0105 p0105 n0105 p0106 n0106 0 tlump
xseg0106 p0106 n0106 p0107 n0107 0 tlump
xseg0107 p0107 n0107 p0108 n0108 0 tlump
xseg0108 p0108 n0108 p0109 n0109 0 tlump
xseg0109 p0109 n0109 p0110 n0110 0 tlump
xseg0110 p0110 n0110 p0111 n0111 0 tlump
xseg0111 p0111 n0111 p0112 n0112 0 tlump
xseg0112 p0112 n0112 p0113 n0113 0 tlump
xseg0113 p0113 n0113 p0114 n0114 0 tlump
xseg0114 p0114 n0114 p0115 n0115 0 tlump
xseg0115 p0115 n0115 p0116 n0116 0 tlump
xseg0116 p0116 n0116 p0117 n0117 0 tlump
xseg0117 p0117 n0117 p0118 n0118 0 tlump
xseg0118 p0118 n0118 p0119 n0119 0 tlump
xseg0119 p0119 n0119 p0120 n0120 0 tlump
xseg0120 p0120 n0120 p0121 n0121 0 tlump
xseg0121 p0121 n0121 p0122 n0122 0 tlump
xseg0122 p0122 n0122 p0123 n0123 0 tlump
xseg0123 p0123 n0123 p0124 n0124 0 tlump
xseg0124 p0124 n0124 p0125 n0125 0 tlump
xseg0125 p0125 n0125 p0126 n0126 0 tlump
xseg0126 p0126 n0126 p0127 n0127 0 tlump
xseg0127 p0127 n0127 p0128 n0128 0 tlump
xseg0128 p0128 n0128 p0129 n0129 0 tlump
xseg0129 p0129 n0129 p0130 n0130 0 tlump
xseg0130 p0130 n0130 p0131 n0131 0 tlump
xseg0131 p0131 n0131 p0132 n0132 0 tlump
xseg0132 p0132 n0132 p0133 n0133 0 tlump
xseg0133 p0133 n0133 p0134 n0134 0 tlump
xseg0134 p0134 n0134 p0135 n0135 0 tlump
xseg0135 p0135 n0135 p0136 n0136 0 tlump
xseg0136 p0136 n0136 p0137 n0137 0 tlump
xseg0137 p0137 n0137 p0138 n0138 0 tlump
xseg0138 p0138 n0138 p0139 n0139 0 tlump
xseg0139 p0139 n0139 p0140 n0140 0 tlump
xseg0140 p0140 n0140 p0141 n0141 0 tlump
xseg0141 p0141 n0141 p0142 n0142 0 tlump
xseg0142 p0142 n0142 p0143 n0143 0 tlump
xseg0143 p0143 n0143 p0144 n0144 0 tlump
xseg0144 p0144 n0144 p0145 n0145 0 tlump
xseg0145 p0145 n0145 p0146 n0146 0 tlump
xseg0146 p0146 n0146 p0147 n0147 0 tlump
xseg0147 p0147 n0147 p0148 n0148 0 tlump
xseg0148 p0148 n0148 p0149 n0149 0 tlump
xseg0149 p0149 n0149 p0150 n0150 0 tlump
xseg0150 p0150 n0150 p0151 n0151 0 tlump
xseg0151 p0151 n0151 p0152 n0152 0 tlump
xseg0152 p0152 n0152 p0153 n0153 0 tlump
xseg0153 p0153 n0153 p0154 n0154 0 tlump
xseg0154 p0154 n0154 p0155 n0155 0 tlump
xseg0155 p0155 n0155 p0156 n0156 0 tlump
xseg0156 p0156 n0156 p0157 n0157 0 tlump
xseg0157 p0157 n0157 p0158 n0158 0 tlump
xseg0158 p0158 n0158 p0159 n0159 0 tlump
xseg0159 p0159 n0159 p0160 n0160 0 tlump
xseg0160 p0160 n0160 p0161 n0161 0 tlump
xseg0161 p0161 n0161 p0162 n0162 0 tlump
xseg0162 p0162 n0162 p0163 n0163 0 tlump
xseg0163 p0163 n0163 p0164 n0164 0 tlump
xseg0164 p0164 n0164 p0165 n0165 0 tlump
xseg0165 p0165 n0165 p0166 n0166 0 tlump
xseg0166 p0166 n0166 p0167 n0167 0 tlump
xseg0167 p0167 n0167 p0168 n0168 0 tlump
xseg0168 p0168 n0168 p0169 n0169 0 tlump
xseg0169 p0169 n0169 p0170 n0170 0 tlump
xseg0170 p0170 n0170 p0171 n0171 0 tlump
xseg0171 p0171 n0171 p0172 n0172 0 tlump
xseg0172 p0172 n0172 p0173 n0173 0 tlump
xseg0173 p0173 n0173 p0174 n0174 0 tlump
xseg0174 p0174 n0174 p0175 n0175 0 tlump
xseg0175 p0175 n0175 p0176 n0176 0 tlump
xseg0176 p0176 n0176 p0177 n0177 0 tlump
xseg0177 p0177 n0177 p0178 n0178 0 tlump
xseg0178 p0178 n0178 p0179 n0179 0 tlump
xseg0179 p0179 n0179 p0180 n0180 0 tlump
xseg0180 p0180 n0180 p0181 n0181 0 tlump
xseg0181 p0181 n0181 p0182 n0182 0 tlump
xseg0182 p0182 n0182 p0183 n0183 0 tlump
xseg0183 p0183 n0183 p0184 n0184 0 tlump
xseg0184 p0184 n0184 p0185 n0185 0 tlump
xseg0185 p0185 n0185 p0186 n0186 0 tlump
xseg0186 p0186 n0186 p0187 n0187 0 tlump
xseg0187 p0187 n0187 p0188 n0188 0 tlump
xseg0188 p0188 n0188 p0189 n0189 0 tlump
xseg0189 p0189 n0189 p0190 n0190 0 tlump
xseg0190 p0190 n0190 p0191 n0191 0 tlump
xseg0191 p0191 n0191 p0192 n0192 0 tlump
xseg0192 p0192 n0192 p0193 n0193 0 tlump
xseg0193 p0193 n0193 p0194 n0194 0 tlump
xseg0194 p0194 n0194 p0195 n0195 0 tlump
xseg0195 p0195 n0195 p0196 n0196 0 tlump
xseg0196 p0196 n0196 p0197 n0197 0 tlump
xseg0197 p0197 n0197 p0198 n0198 0 tlump
xseg0198 p0198 n0198 p0199 n0199 0 tlump
xseg0199 p0199 n0199 p0200 n0200 0 tlump
xseg0200 p0200 n0200 p0201 n0201 0 tlump
xseg0201 p0201 n0201 p0202 n0202 0 tlump
xseg0202 p0202 n0202 p0203 n0203 0 tlump
xseg0203 p0203 n0203 p0204 n0204 0 tlump
xseg0204 p0204 n0204 p0205 n0205 0 tlump
xseg0205 p0205 n0205 p0206 n0206 0 tlump
xseg0206 p0206 n0206 p0207 n0207 0 tlump
xseg0207 p0207 n0207 p0208 n0208 0 tlump
xseg0208 p0208 n0208 p0209 n0209 0 tlump
xseg0209 p0209 n0209 p0210 n0210 0 tlump
xseg0210 p0210 n0210 p0211 n0211 0 tlump
xseg0211 p0211 n0211 p0212 n0212 0 tlump
xseg0212 p0212 n0212 p0213 n0213 0 tlump
xseg0213 p0213 n0213 p0214 n0214 0 tlump
xseg0214 p0214 n0214 p0215 n0215 0 tlump
xseg0215 p0215 n0215 p0216 n0216 0 tlump
xseg0216 p0216 n0216 p0217 n0217 0 tlump
xseg0217 p0217 n0217 p0218 n0218 0 tlump
xseg0218 p0218 n0218 p0219 n0219 0 tlump
xseg0219 p0219 n0219 p0220 n0220 0 tlump
xseg0220 p0220 n0220 p0221 n0221 0 tlump
xseg0221 p0221 n0221 p0222 n0222 0 tlump
xseg0222 p0222 n0222 p0223 n0223 0 tlump
xseg0223 p0223 n0223 p0224 n0224 0 tlump
xseg0224 p0224 n0224 p0225 n0225 0 tlump
xseg0225 p0225 n0225 p0226 n0226 0 tlump
xseg0226 p0226 n0226 p0227 n0227 0 tlump
xseg0227 p0227 n0227 p0228 n0228 0 tlump
xseg0228 p0228 n0228 p0229 n0229 0 tlump
xseg0229 p0229 n0229 p0230 n0230 0 tlump
xseg0230 p0230 n0230 p0231 n0231 0 tlump
xseg0231 p0231 n0231 p0232 n0232 0 tlump
xseg0232 p0232 n0232 p0233 n0233 0 tlump
xseg0233 p0233 n0233 p0234 n0234 0 tlump
xseg0234 p0234 n0234 p0235 n0235 0 tlump
xseg0235 p0235 n0235 p0236 n0236 0 tlump
xseg0236 p0236 n0236 p0237 n0237 0 tlump
xseg0237 p0237 n0237 p0238 n0238 0 tlump
xseg0238 p0238 n0238 p0239 n0239 0 tlump
xseg0239 p0239 n0239 p0240 n0240 0 tlump
xseg0240 p0240 n0240 p0241 n0241 0 tlump
xseg0241 p0241 n0241 p0242 n0242 0 tlump
xseg0242 p0242 n0242 p0243 n0243 0 tlump
xseg0243 p0243 n0243 p0244 n0244 0 tlump
xseg0244 p0244 n0244 p0245 n0245 0 tlump
xseg0245 p0245 n0245 p0246 n0246 0 tlump
xseg0246 p0246 n0246 p0247 n0247 0 tlump
xseg0247 p0247 n0247 p0248 n0248 0 tlump
xseg0248 p0248 n0248 p0249 n0249 0 tlump
xseg0249 p0249 n0249 p0250 n0250 0 tlump
xseg0250 p0250 n0250 p0251 n0251 0 tlump
xseg0251 p0251 n0251 p0252 n0252 0 tlump
xseg0252 p0252 n0252 p0253 n0253 0 tlump
xseg0253 p0253 n0253 p0254 n0254 0 tlump
xseg0254 p0254 n0254 p0255 n0255 0 tlump
xseg0255 p0255 n0255 p0256 n0256 0 tlump
xseg0256 p0256 n0256 p0257 n0257 0 tlump
xseg0257 p0257 n0257 p0258 n0258 0 tlump
xseg0258 p0258 n0258 p0259 n0259 0 tlump
xseg0259 p0259 n0259 p0260 n0260 0 tlump
xseg0260 p0260 n0260 p0261 n0261 0 tlump
xseg0261 p0261 n0261 p0262 n0262 0 tlump
xseg0262 p0262 n0262 p0263 n0263 0 tlump
xseg0263 p0263 n0263 p0264 n0264 0 tlump
xseg0264 p0264 n0264 p0265 n0265 0 tlump
xseg0265 p0265 n0265 p0266 n0266 0 tlump
xseg0266 p0266 n0266 p0267 n0267 0 tlump
xseg0267 p0267 n0267 p0268 n0268 0 tlump
xseg0268 p0268 n0268 p0269 n0269 0 tlump
xseg0269 p0269 n0269 p0270 n0270 0 tlump
xseg0270 p0270 n0270 p0271 n0271 0 tlump
xseg0271 p0271 n0271 p0272 n0272 0 tlump
xseg0272 p0272 n0272 p0273 n0273 0 tlump
xseg0273 p0273 n0273 p0274 n0274 0 tlump
xseg0274 p0274 n0274 p0275 n0275 0 tlump
xseg0275 p0275 n0275 p0276 n0276 0 tlump
xseg0276 p0276 n0276 p0277 n0277 0 tlump
xseg0277 p0277 n0277 p0278 n0278 0 tlump
xseg0278 p0278 n0278 p0279 n0279 0 tlump
xseg0279 p0279 n0279 p0280 n0280 0 tlump
xseg0280 p0280 n0280 p0281 n0281 0 tlump
xseg0281 p0281 n0281 p0282 n0282 0 tlump
xseg0282 p0282 n0282 p0283 n0283 0 tlump
xseg0283 p0283 n0283 p0284 n0284 0 tlump
xseg0284 p0284 n0284 p0285 n0285 0 tlump
xseg0285 p0285 n0285 p0286 n0286 0 tlump
xseg0286 p0286 n0286 p0287 n0287 0 tlump
xseg0287 p0287 n0287 p0288 n0288 0 tlump
xseg0288 p0288 n0288 p0289 n0289 0 tlump
xseg0289 p0289 n0289 p0290 n0290 0 tlump
xseg0290 p0290 n0290 p0291 n0291 0 tlump
xseg0291 p0291 n0291 p0292 n0292 0 tlump
xseg0292 p0292 n0292 p0293 n0293 0 tlump
xseg0293 p0293 n0293 p0294 n0294 0 tlump
xseg0294 p0294 n0294 p0295 n0295 0 tlump
xseg0295 p0295 n0295 p0296 n0296 0 tlump
xseg0296 p0296 n0296 p0297 n0297 0 tlump
xseg0297 p0297 n0297 p0298 n0298 0 tlump
xseg0298 p0298 n0298 p0299 n0299 0 tlump
xseg0299 p0299 n0299 p0300 n0300 0 tlump
xseg0300 p0300 n0300 p0301 n0301 0 tlump
xseg0301 p0301 n0301 p0302 n0302 0 tlump
xseg0302 p0302 n0302 p0303 n0303 0 tlump
xseg0303 p0303 n0303 p0304 n0304 0 tlump
xseg0304 p0304 n0304 p0305 n0305 0 tlump
xseg0305 p0305 n0305 p0306 n0306 0 tlump
xseg0306 p0306 n0306 p0307 n0307 0 tlump
xseg0307 p0307 n0307 p0308 n0308 0 tlump
xseg0308 p0308 n0308 p0309 n0309 0 tlump
xseg0309 p0309 n0309 p0310 n0310 0 tlump
xseg0310 p0310 n0310 p0311 n0311 0 tlump
xseg0311 p0311 n0311 p0312 n0312 0 tlump
xseg0312 p0312 n0312 p0313 n0313 0 tlump
xseg0313 p0313 n0313 p0314 n0314 0 tlump
xseg0314 p0314 n0314 p0315 n0315 0 tlump
xseg0315 p0315 n0315 p0316 n0316 0 tlump
xseg0316 p0316 n0316 p0317 n0317 0 tlump
xseg0317 p0317 n0317 p0318 n0318 0 tlump
xseg0318 p0318 n0318 p0319 n0319 0 tlump
xseg0319 p0319 n0319 p0320 n0320 0 tlump
xseg0320 p0320 n0320 p0321 n0321 0 tlump
xseg0321 p0321 n0321 p0322 n0322 0 tlump
xseg0322 p0322 n0322 p0323 n0323 0 tlump
xseg0323 p0323 n0323 p0324 n0324 0 tlump
xseg0324 p0324 n0324 p0325 n0325 0 tlump
xseg0325 p0325 n0325 p0326 n0326 0 tlump
xseg0326 p0326 n0326 p0327 n0327 0 tlump
xseg0327 p0327 n0327 p0328 n0328 0 tlump
xseg0328 p0328 n0328 p0329 n0329 0 tlump
xseg0329 p0329 n0329 p0330 n0330 0 tlump
xseg0330 p0330 n0330 p0331 n0331 0 tlump
xseg0331 p0331 n0331 p0332 n0332 0 tlump
xseg0332 p0332 n0332 p0333 n0333 0 tlump
xseg0333 p0333 n0333 p0334 n0334 0 tlump
xseg0334 p0334 n0334 p0335 n0335 0 tlump
xseg0335 p0335 n0335 p0336 n0336 0 tlump
xseg0336 p0336 n0336 p0337 n0337 0 tlump
xseg0337 p0337 n0337 p0338 n0338 0 tlump
xseg0338 p0338 n0338 p0339 n0339 0 tlump
xseg0339 p0339 n0339 p0340 n0340 0 tlump
xseg0340 p0340 n0340 p0341 n0341 0 tlump
xseg0341 p0341 n0341 p0342 n0342 0 tlump
xseg0342 p0342 n0342 p0343 n0343 0 tlump
xseg0343 p0343 n0343 p0344 n0344 0 tlump
xseg0344 p0344 n0344 p0345 n0345 0 tlump
xseg0345 p0345 n0345 p0346 n0346 0 tlump
xseg0346 p0346 n0346 p0347 n0347 0 tlump
xseg0347 p0347 n0347 p0348 n0348 0 tlump
xseg0348 p0348 n0348 p0349 n0349 0 tlump
xseg0349 p0349 n0349 p0350 n0350 0 tlump
xseg0350 p0350 n0350 p0351 n0351 0 tlump
xseg0351 p0351 n0351 p0352 n0352 0 tlump
xseg0352 p0352 n0352 p0353 n0353 0 tlump
xseg0353 p0353 n0353 p0354 n0354 0 tlump
xseg0354 p0354 n0354 p0355 n0355 0 tlump
xseg0355 p0355 n0355 p0356 n0356 0 tlump
xseg0356 p0356 n0356 p0357 n0357 0 tlump
xseg0357 p0357 n0357 p0358 n0358 0 tlump
xseg0358 p0358 n0358 p0359 n0359 0 tlump
xseg0359 p0359 n0359 p0360 n0360 0 tlump
xseg0360 p0360 n0360 p0361 n0361 0 tlump
xseg0361 p0361 n0361 p0362 n0362 0 tlump
xseg0362 p0362 n0362 p0363 n0363 0 tlump
xseg0363 p0363 n0363 p0364 n0364 0 tlump
xseg0364 p0364 n0364 p0365 n0365 0 tlump
xseg0365 p0365 n0365 p0366 n0366 0 tlump
xseg0366 p0366 n0366 p0367 n0367 0 tlump
xseg0367 p0367 n0367 p0368 n0368 0 tlump
xseg0368 p0368 n0368 p0369 n0369 0 tlump
xseg0369 p0369 n0369 p0370 n0370 0 tlump
xseg0370 p0370 n0370 p0371 n0371 0 tlump
xseg0371 p0371 n0371 p0372 n0372 0 tlump
xseg0372 p0372 n0372 p0373 n0373 0 tlump
xseg0373 p0373 n0373 p0374 n0374 0 tlump
xseg0374 p0374 n0374 p0375 n0375 0 tlump
xseg0375 p0375 n0375 p0376 n0376 0 tlump
xseg0376 p0376 n0376 p0377 n0377 0 tlump
xseg0377 p0377 n0377 p0378 n0378 0 tlump
xseg0378 p0378 n0378 p0379 n0379 0 tlump
xseg0379 p0379 n0379 p0380 n0380 0 tlump
xseg0380 p0380 n0380 p0381 n0381 0 tlump
xseg0381 p0381 n0381 p0382 n0382 0 tlump
xseg0382 p0382 n0382 p0383 n0383 0 tlump
xseg0383 p0383 n0383 p0384 n0384 0 tlump
xseg0384 p0384 n0384 p0385 n0385 0 tlump
xseg0385 p0385 n0385 p0386 n0386 0 tlump
xseg0386 p0386 n0386 p0387 n0387 0 tlump
xseg0387 p0387 n0387 p0388 n0388 0 tlump
xseg0388 p0388 n0388 p0389 n0389 0 tlump
xseg0389 p0389 n0389 p0390 n0390 0 tlump
xseg0390 p0390 n0390 p0391 n0391 0 tlump
xseg0391 p0391 n0391 p0392 n0392 0 tlump
xseg0392 p0392 n0392 p0393 n0393 0 tlump
xseg0393 p0393 n0393 p0394 n0394 0 tlump
xseg0394 p0394 n0394 p0395 n0395 0 tlump
xseg0395 p0395 n0395 p0396 n0396 0 tlump
xseg0396 p0396 n0396 p0397 n0397 0 tlump
xseg0397 p0397 n0397 p0398 n0398 0 tlump
xseg0398 p0398 n0398 p0399 n0399 0 tlump
xseg0399 p0399 n0399 p0400 n0400 0 tlump
xseg0400 p0400 n0400 p0401 n0401 0 tlump
xseg0401 p0401 n0401 p0402 n0402 0 tlump
xseg0402 p0402 n0402 p0403 n0403 0 tlump
xseg0403 p0403 n0403 p0404 n0404 0 tlump
xseg0404 p0404 n0404 p0405 n0405 0 tlump
xseg0405 p0405 n0405 p0406 n0406 0 tlump
xseg0406 p0406 n0406 p0407 n0407 0 tlump
xseg0407 p0407 n0407 p0408 n0408 0 tlump
xseg0408 p0408 n0408 p0409 n0409 0 tlump
xseg0409 p0409 n0409 p0410 n0410 0 tlump
xseg0410 p0410 n0410 p0411 n0411 0 tlump
xseg0411 p0411 n0411 p0412 n0412 0 tlump
xseg0412 p0412 n0412 p0413 n0413 0 tlump
xseg0413 p0413 n0413 p0414 n0414 0 tlump
xseg0414 p0414 n0414 p0415 n0415 0 tlump
xseg0415 p0415 n0415 p0416 n0416 0 tlump
xseg0416 p0416 n0416 p0417 n0417 0 tlump
xseg0417 p0417 n0417 p0418 n0418 0 tlump
xseg0418 p0418 n0418 p0419 n0419 0 tlump
xseg0419 p0419 n0419 p0420 n0420 0 tlump
xseg0420 p0420 n0420 p0421 n0421 0 tlump
xseg0421 p0421 n0421 p0422 n0422 0 tlump
xseg0422 p0422 n0422 p0423 n0423 0 tlump
xseg0423 p0423 n0423 p0424 n0424 0 tlump
xseg0424 p0424 n0424 p0425 n0425 0 tlump
xseg0425 p0425 n0425 p0426 n0426 0 tlump
xseg0426 p0426 n0426 p0427 n0427 0 tlump
xseg0427 p0427 n0427 p0428 n0428 0 tlump
xseg0428 p0428 n0428 p0429 n0429 0 tlump
xseg0429 p0429 n0429 p0430 n0430 0 tlump
xseg0430 p0430 n0430 p0431 n0431 0 tlump
xseg0431 p0431 n0431 p0432 n0432 0 tlump
xseg0432 p0432 n0432 p0433 n0433 0 tlump
xseg0433 p0433 n0433 p0434 n0434 0 tlump
xseg0434 p0434 n0434 p0435 n0435 0 tlump
xseg0435 p0435 n0435 p0436 n0436 0 tlump
xseg0436 p0436 n0436 p0437 n0437 0 tlump
xseg0437 p0437 n0437 p0438 n0438 0 tlump
xseg0438 p0438 n0438 p0439 n0439 0 tlump
xseg0439 p0439 n0439 p0440 n0440 0 tlump
xseg0440 p0440 n0440 p0441 n0441 0 tlump
xseg0441 p0441 n0441 p0442 n0442 0 tlump
xseg0442 p0442 n0442 p0443 n0443 0 tlump
xseg0443 p0443 n0443 p0444 n0444 0 tlump
xseg0444 p0444 n0444 p0445 n0445 0 tlump
xseg0445 p0445 n0445 p0446 n0446 0 tlump
xseg0446 p0446 n0446 p0447 n0447 0 tlump
xseg0447 p0447 n0447 p0448 n0448 0 tlump
xseg0448 p0448 n0448 p0449 n0449 0 tlump
xseg0449 p0449 n0449 p0450 n0450 0 tlump
xseg0450 p0450 n0450 p0451 n0451 0 tlump
xseg0451 p0451 n0451 p0452 n0452 0 tlump
xseg0452 p0452 n0452 p0453 n0453 0 tlump
xseg0453 p0453 n0453 p0454 n0454 0 tlump
xseg0454 p0454 n0454 p0455 n0455 0 tlump
xseg0455 p0455 n0455 p0456 n0456 0 tlump
xseg0456 p0456 n0456 p0457 n0457 0 tlump
xseg0457 p0457 n0457 p0458 n0458 0 tlump
xseg0458 p0458 n0458 p0459 n0459 0 tlump
xseg0459 p0459 n0459 p0460 n0460 0 tlump
xseg0460 p0460 n0460 p0461 n0461 0 tlump
xseg0461 p0461 n0461 p0462 n0462 0 tlump
xseg0462 p0462 n0462 p0463 n0463 0 tlump
xseg0463 p0463 n0463 p0464 n0464 0 tlump
xseg0464 p0464 n0464 p0465 n0465 0 tlump
xseg0465 p0465 n0465 p0466 n0466 0 tlump
xseg0466 p0466 n0466 p0467 n0467 0 tlump
xseg0467 p0467 n0467 p0468 n0468 0 tlump
xseg0468 p0468 n0468 p0469 n0469 0 tlump
xseg0469 p0469 n0469 p0470 n0470 0 tlump
xseg0470 p0470 n0470 p0471 n0471 0 tlump
xseg0471 p0471 n0471 p0472 n0472 0 tlump
xseg0472 p0472 n0472 p0473 n0473 0 tlump
xseg0473 p0473 n0473 p0474 n0474 0 tlump
xseg0474 p0474 n0474 p0475 n0475 0 tlump
xseg0475 p0475 n0475 p0476 n0476 0 tlump
xseg0476 p0476 n0476 p0477 n0477 0 tlump
xseg0477 p0477 n0477 p0478 n0478 0 tlump
xseg0478 p0478 n0478 p0479 n0479 0 tlump
xseg0479 p0479 n0479 p0480 n0480 0 tlump
xseg0480 p0480 n0480 p0481 n0481 0 tlump
xseg0481 p0481 n0481 p0482 n0482 0 tlump
xseg0482 p0482 n0482 p0483 n0483 0 tlump
xseg0483 p0483 n0483 p0484 n0484 0 tlump
xseg0484 p0484 n0484 p0485 n0485 0 tlump
xseg0485 p0485 n0485 p0486 n0486 0 tlump
xseg0486 p0486 n0486 p0487 n0487 0 tlump
xseg0487 p0487 n0487 p0488 n0488 0 tlump
xseg0488 p0488 n0488 p0489 n0489 0 tlump
xseg0489 p0489 n0489 p0490 n0490 0 tlump
xseg0490 p0490 n0490 p0491 n0491 0 tlump
xseg0491 p0491 n0491 p0492 n0492 0 tlump
xseg0492 p0492 n0492 p0493 n0493 0 tlump
xseg0493 p0493 n0493 p0494 n0494 0 tlump
xseg0494 p0494 n0494 p0495 n0495 0 tlump
xseg0495 p0495 n0495 p0496 n0496 0 tlump
xseg0496 p0496 n0496 p0497 n0497 0 tlump
xseg0497 p0497 n0497 p0498 n0498 0 tlump
xseg0498 p0498 n0498 p0499 n0499 0 tlump
xseg0499 p0499 n0499 p0500 n0500 0 tlump
xseg0500 p0500 n0500 p0501 n0501 0 tlump
xseg0501 p0501 n0501 p0502 n0502 0 tlump
xseg0502 p0502 n0502 p0503 n0503 0 tlump
xseg0503 p0503 n0503 p0504 n0504 0 tlump
xseg0504 p0504 n0504 p0505 n0505 0 tlump
xseg0505 p0505 n0505 p0506 n0506 0 tlump
xseg0506 p0506 n0506 p0507 n0507 0 tlump
xseg0507 p0507 n0507 p0508 n0508 0 tlump
xseg0508 p0508 n0508 p0509 n0509 0 tlump
xseg0509 p0509 n0509 p0510 n0510 0 tlump
xseg0510 p0510 n0510 p0511 n0511 0 tlump
xseg0511 p0511 n0511 p0512 n0512 0 tlump
xseg0512 p0512 n0512 p0513 n0513 0 tlump
xseg0513 p0513 n0513 p0514 n0514 0 tlump
xseg0514 p0514 n0514 p0515 n0515 0 tlump
xseg0515 p0515 n0515 p0516 n0516 0 tlump
xseg0516 p0516 n0516 p0517 n0517 0 tlump
xseg0517 p0517 n0517 p0518 n0518 0 tlump
xseg0518 p0518 n0518 p0519 n0519 0 tlump
xseg0519 p0519 n0519 p0520 n0520 0 tlump
xseg0520 p0520 n0520 p0521 n0521 0 tlump
xseg0521 p0521 n0521 p0522 n0522 0 tlump
xseg0522 p0522 n0522 p0523 n0523 0 tlump
xseg0523 p0523 n0523 p0524 n0524 0 tlump
xseg0524 p0524 n0524 p0525 n0525 0 tlump
xseg0525 p0525 n0525 p0526 n0526 0 tlump
xseg0526 p0526 n0526 p0527 n0527 0 tlump
xseg0527 p0527 n0527 p0528 n0528 0 tlump
xseg0528 p0528 n0528 p0529 n0529 0 tlump
xseg0529 p0529 n0529 p0530 n0530 0 tlump
xseg0530 p0530 n0530 p0531 n0531 0 tlump
xseg0531 p0531 n0531 p0532 n0532 0 tlump
xseg0532 p0532 n0532 p0533 n0533 0 tlump
xseg0533 p0533 n0533 p0534 n0534 0 tlump
xseg0534 p0534 n0534 p0535 n0535 0 tlump
xseg0535 p0535 n0535 p0536 n0536 0 tlump
xseg0536 p0536 n0536 p0537 n0537 0 tlump
xseg0537 p0537 n0537 p0538 n0538 0 tlump
xseg0538 p0538 n0538 p0539 n0539 0 tlump
xseg0539 p0539 n0539 p0540 n0540 0 tlump
xseg0540 p0540 n0540 p0541 n0541 0 tlump
xseg0541 p0541 n0541 p0542 n0542 0 tlump
xseg0542 p0542 n0542 p0543 n0543 0 tlump
xseg0543 p0543 n0543 p0544 n0544 0 tlump
xseg0544 p0544 n0544 p0545 n0545 0 tlump
xseg0545 p0545 n0545 p0546 n0546 0 tlump
xseg0546 p0546 n0546 p0547 n0547 0 tlump
xseg0547 p0547 n0547 p0548 n0548 0 tlump
xseg0548 p0548 n0548 p0549 n0549 0 tlump
xseg0549 p0549 n0549 p0550 n0550 0 tlump
xseg0550 p0550 n0550 p0551 n0551 0 tlump
xseg0551 p0551 n0551 p0552 n0552 0 tlump
xseg0552 p0552 n0552 p0553 n0553 0 tlump
xseg0553 p0553 n0553 p0554 n0554 0 tlump
xseg0554 p0554 n0554 p0555 n0555 0 tlump
xseg0555 p0555 n0555 p0556 n0556 0 tlump
xseg0556 p0556 n0556 p0557 n0557 0 tlump
xseg0557 p0557 n0557 p0558 n0558 0 tlump
xseg0558 p0558 n0558 p0559 n0559 0 tlump
xseg0559 p0559 n0559 p0560 n0560 0 tlump
xseg0560 p0560 n0560 p0561 n0561 0 tlump
xseg0561 p0561 n0561 p0562 n0562 0 tlump
xseg0562 p0562 n0562 p0563 n0563 0 tlump
xseg0563 p0563 n0563 p0564 n0564 0 tlump
xseg0564 p0564 n0564 p0565 n0565 0 tlump
xseg0565 p0565 n0565 p0566 n0566 0 tlump
xseg0566 p0566 n0566 p0567 n0567 0 tlump
xseg0567 p0567 n0567 p0568 n0568 0 tlump
xseg0568 p0568 n0568 p0569 n0569 0 tlump
xseg0569 p0569 n0569 p0570 n0570 0 tlump
xseg0570 p0570 n0570 p0571 n0571 0 tlump
xseg0571 p0571 n0571 p0572 n0572 0 tlump
xseg0572 p0572 n0572 p0573 n0573 0 tlump
xseg0573 p0573 n0573 p0574 n0574 0 tlump
xseg0574 p0574 n0574 p0575 n0575 0 tlump
xseg0575 p0575 n0575 p0576 n0576 0 tlump
xseg0576 p0576 n0576 p0577 n0577 0 tlump
xseg0577 p0577 n0577 p0578 n0578 0 tlump
xseg0578 p0578 n0578 p0579 n0579 0 tlump
xseg0579 p0579 n0579 p0580 n0580 0 tlump
xseg0580 p0580 n0580 p0581 n0581 0 tlump
xseg0581 p0581 n0581 p0582 n0582 0 tlump
xseg0582 p0582 n0582 p0583 n0583 0 tlump
xseg0583 p0583 n0583 p0584 n0584 0 tlump
xseg0584 p0584 n0584 p0585 n0585 0 tlump
xseg0585 p0585 n0585 p0586 n0586 0 tlump
xseg0586 p0586 n0586 p0587 n0587 0 tlump
xseg0587 p0587 n0587 p0588 n0588 0 tlump
xseg0588 p0588 n0588 p0589 n0589 0 tlump
xseg0589 p0589 n0589 p0590 n0590 0 tlump
xseg0590 p0590 n0590 p0591 n0591 0 tlump
xseg0591 p0591 n0591 p0592 n0592 0 tlump
xseg0592 p0592 n0592 p0593 n0593 0 tlump
xseg0593 p0593 n0593 p0594 n0594 0 tlump
xseg0594 p0594 n0594 p0595 n0595 0 tlump
xseg0595 p0595 n0595 p0596 n0596 0 tlump
xseg0596 p0596 n0596 p0597 n0597 0 tlump
xseg0597 p0597 n0597 p0598 n0598 0 tlump
xseg0598 p0598 n0598 p0599 n0599 0 tlump
xseg0599 p0599 n0599 p0600 n0600 0 tlump
xseg0600 p0600 n0600 p0601 n0601 0 tlump
xseg0601 p0601 n0601 p0602 n0602 0 tlump
xseg0602 p0602 n0602 p0603 n0603 0 tlump
xseg0603 p0603 n0603 p0604 n0604 0 tlump
xseg0604 p0604 n0604 p0605 n0605 0 tlump
xseg0605 p0605 n0605 p0606 n0606 0 tlump
xseg0606 p0606 n0606 p0607 n0607 0 tlump
xseg0607 p0607 n0607 p0608 n0608 0 tlump
xseg0608 p0608 n0608 p0609 n0609 0 tlump
xseg0609 p0609 n0609 p0610 n0610 0 tlump
xseg0610 p0610 n0610 p0611 n0611 0 tlump
xseg0611 p0611 n0611 p0612 n0612 0 tlump
xseg0612 p0612 n0612 p0613 n0613 0 tlump
xseg0613 p0613 n0613 p0614 n0614 0 tlump
xseg0614 p0614 n0614 p0615 n0615 0 tlump
xseg0615 p0615 n0615 p0616 n0616 0 tlump
xseg0616 p0616 n0616 p0617 n0617 0 tlump
xseg0617 p0617 n0617 p0618 n0618 0 tlump
xseg0618 p0618 n0618 p0619 n0619 0 tlump
xseg0619 p0619 n0619 p0620 n0620 0 tlump
xseg0620 p0620 n0620 p0621 n0621 0 tlump
xseg0621 p0621 n0621 p0622 n0622 0 tlump
xseg0622 p0622 n0622 p0623 n0623 0 tlump
xseg0623 p0623 n0623 p0624 n0624 0 tlump
xseg0624 p0624 n0624 p0625 n0625 0 tlump
xseg0625 p0625 n0625 p0626 n0626 0 tlump
xseg0626 p0626 n0626 p0627 n0627 0 tlump
xseg0627 p0627 n0627 p0628 n0628 0 tlump
xseg0628 p0628 n0628 p0629 n0629 0 tlump
xseg0629 p0629 n0629 p0630 n0630 0 tlump
xseg0630 p0630 n0630 p0631 n0631 0 tlump
xseg0631 p0631 n0631 p0632 n0632 0 tlump
xseg0632 p0632 n0632 p0633 n0633 0 tlump
xseg0633 p0633 n0633 p0634 n0634 0 tlump
xseg0634 p0634 n0634 p0635 n0635 0 tlump
xseg0635 p0635 n0635 p0636 n0636 0 tlump
xseg0636 p0636 n0636 p0637 n0637 0 tlump
xseg0637 p0637 n0637 p0638 n0638 0 tlump
xseg0638 p0638 n0638 p0639 n0639 0 tlump
xseg0639 p0639 n0639 p0640 n0640 0 tlump
xseg0640 p0640 n0640 p0641 n0641 0 tlump
xseg0641 p0641 n0641 p0642 n0642 0 tlump
xseg0642 p0642 n0642 p0643 n0643 0 tlump
xseg0643 p0643 n0643 p0644 n0644 0 tlump
xseg0644 p0644 n0644 p0645 n0645 0 tlump
xseg0645 p0645 n0645 p0646 n0646 0 tlump
xseg0646 p0646 n0646 p0647 n0647 0 tlump
xseg0647 p0647 n0647 p0648 n0648 0 tlump
xseg0648 p0648 n0648 p0649 n0649 0 tlump
xseg0649 p0649 n0649 p0650 n0650 0 tlump
xseg0650 p0650 n0650 p0651 n0651 0 tlump
xseg0651 p0651 n0651 p0652 n0652 0 tlump
xseg0652 p0652 n0652 p0653 n0653 0 tlump
xseg0653 p0653 n0653 p0654 n0654 0 tlump
xseg0654 p0654 n0654 p0655 n0655 0 tlump
xseg0655 p0655 n0655 p0656 n0656 0 tlump
xseg0656 p0656 n0656 p0657 n0657 0 tlump
xseg0657 p0657 n0657 p0658 n0658 0 tlump
xseg0658 p0658 n0658 p0659 n0659 0 tlump
xseg0659 p0659 n0659 p0660 n0660 0 tlump
xseg0660 p0660 n0660 p0661 n0661 0 tlump
xseg0661 p0661 n0661 p0662 n0662 0 tlump
xseg0662 p0662 n0662 p0663 n0663 0 tlump
xseg0663 p0663 n0663 p0664 n0664 0 tlump
xseg0664 p0664 n0664 p0665 n0665 0 tlump
xseg0665 p0665 n0665 p0666 n0666 0 tlump
xseg0666 p0666 n0666 p0667 n0667 0 tlump
xseg0667 p0667 n0667 p0668 n0668 0 tlump
xseg0668 p0668 n0668 p0669 n0669 0 tlump
xseg0669 p0669 n0669 p0670 n0670 0 tlump
xseg0670 p0670 n0670 p0671 n0671 0 tlump
xseg0671 p0671 n0671 p0672 n0672 0 tlump
xseg0672 p0672 n0672 p0673 n0673 0 tlump
xseg0673 p0673 n0673 p0674 n0674 0 tlump
xseg0674 p0674 n0674 p0675 n0675 0 tlump
xseg0675 p0675 n0675 p0676 n0676 0 tlump
xseg0676 p0676 n0676 p0677 n0677 0 tlump
xseg0677 p0677 n0677 p0678 n0678 0 tlump
xseg0678 p0678 n0678 p0679 n0679 0 tlump
xseg0679 p0679 n0679 p0680 n0680 0 tlump
xseg0680 p0680 n0680 p0681 n0681 0 tlump
xseg0681 p0681 n0681 p0682 n0682 0 tlump
xseg0682 p0682 n0682 p0683 n0683 0 tlump
xseg0683 p0683 n0683 p0684 n0684 0 tlump
xseg0684 p0684 n0684 p0685 n0685 0 tlump
xseg0685 p0685 n0685 p0686 n0686 0 tlump
xseg0686 p0686 n0686 p0687 n0687 0 tlump
xseg0687 p0687 n0687 p0688 n0688 0 tlump
xseg0688 p0688 n0688 p0689 n0689 0 tlump
xseg0689 p0689 n0689 p0690 n0690 0 tlump
xseg0690 p0690 n0690 p0691 n0691 0 tlump
xseg0691 p0691 n0691 p0692 n0692 0 tlump
xseg0692 p0692 n0692 p0693 n0693 0 tlump
xseg0693 p0693 n0693 p0694 n0694 0 tlump
xseg0694 p0694 n0694 p0695 n0695 0 tlump
xseg0695 p0695 n0695 p0696 n0696 0 tlump
xseg0696 p0696 n0696 p0697 n0697 0 tlump
xseg0697 p0697 n0697 p0698 n0698 0 tlump
xseg0698 p0698 n0698 p0699 n0699 0 tlump
xseg0699 p0699 n0699 p0700 n0700 0 tlump
xseg0700 p0700 n0700 p0701 n0701 0 tlump
xseg0701 p0701 n0701 p0702 n0702 0 tlump
xseg0702 p0702 n0702 p0703 n0703 0 tlump
xseg0703 p0703 n0703 p0704 n0704 0 tlump
xseg0704 p0704 n0704 p0705 n0705 0 tlump
xseg0705 p0705 n0705 p0706 n0706 0 tlump
xseg0706 p0706 n0706 p0707 n0707 0 tlump
xseg0707 p0707 n0707 p0708 n0708 0 tlump
xseg0708 p0708 n0708 p0709 n0709 0 tlump
xseg0709 p0709 n0709 p0710 n0710 0 tlump
xseg0710 p0710 n0710 p0711 n0711 0 tlump
xseg0711 p0711 n0711 p0712 n0712 0 tlump
xseg0712 p0712 n0712 p0713 n0713 0 tlump
xseg0713 p0713 n0713 p0714 n0714 0 tlump
xseg0714 p0714 n0714 p0715 n0715 0 tlump
xseg0715 p0715 n0715 p0716 n0716 0 tlump
xseg0716 p0716 n0716 p0717 n0717 0 tlump
xseg0717 p0717 n0717 p0718 n0718 0 tlump
xseg0718 p0718 n0718 p0719 n0719 0 tlump
xseg0719 p0719 n0719 p0720 n0720 0 tlump
xseg0720 p0720 n0720 p0721 n0721 0 tlump
xseg0721 p0721 n0721 p0722 n0722 0 tlump
xseg0722 p0722 n0722 p0723 n0723 0 tlump
xseg0723 p0723 n0723 p0724 n0724 0 tlump
xseg0724 p0724 n0724 p0725 n0725 0 tlump
xseg0725 p0725 n0725 p0726 n0726 0 tlump
xseg0726 p0726 n0726 p0727 n0727 0 tlump
xseg0727 p0727 n0727 p0728 n0728 0 tlump
xseg0728 p0728 n0728 p0729 n0729 0 tlump
xseg0729 p0729 n0729 p0730 n0730 0 tlump
xseg0730 p0730 n0730 p0731 n0731 0 tlump
xseg0731 p0731 n0731 p0732 n0732 0 tlump
xseg0732 p0732 n0732 p0733 n0733 0 tlump
xseg0733 p0733 n0733 p0734 n0734 0 tlump
xseg0734 p0734 n0734 p0735 n0735 0 tlump
xseg0735 p0735 n0735 p0736 n0736 0 tlump
xseg0736 p0736 n0736 p0737 n0737 0 tlump
xseg0737 p0737 n0737 p0738 n0738 0 tlump
xseg0738 p0738 n0738 p0739 n0739 0 tlump
xseg0739 p0739 n0739 p0740 n0740 0 tlump
xseg0740 p0740 n0740 p0741 n0741 0 tlump
xseg0741 p0741 n0741 p0742 n0742 0 tlump
xseg0742 p0742 n0742 p0743 n0743 0 tlump
xseg0743 p0743 n0743 p0744 n0744 0 tlump
xseg0744 p0744 n0744 p0745 n0745 0 tlump
xseg0745 p0745 n0745 p0746 n0746 0 tlump
xseg0746 p0746 n0746 p0747 n0747 0 tlump
xseg0747 p0747 n0747 p0748 n0748 0 tlump
xseg0748 p0748 n0748 p0749 n0749 0 tlump
xseg0749 p0749 n0749 p0750 n0750 0 tlump
xseg0750 p0750 n0750 p0751 n0751 0 tlump
xseg0751 p0751 n0751 p0752 n0752 0 tlump
xseg0752 p0752 n0752 p0753 n0753 0 tlump
xseg0753 p0753 n0753 p0754 n0754 0 tlump
xseg0754 p0754 n0754 p0755 n0755 0 tlump
xseg0755 p0755 n0755 p0756 n0756 0 tlump
xseg0756 p0756 n0756 p0757 n0757 0 tlump
xseg0757 p0757 n0757 p0758 n0758 0 tlump
xseg0758 p0758 n0758 p0759 n0759 0 tlump
xseg0759 p0759 n0759 p0760 n0760 0 tlump
xseg0760 p0760 n0760 p0761 n0761 0 tlump
xseg0761 p0761 n0761 p0762 n0762 0 tlump
xseg0762 p0762 n0762 p0763 n0763 0 tlump
xseg0763 p0763 n0763 p0764 n0764 0 tlump
xseg0764 p0764 n0764 p0765 n0765 0 tlump
xseg0765 p0765 n0765 p0766 n0766 0 tlump
xseg0766 p0766 n0766 p0767 n0767 0 tlump
xseg0767 p0767 n0767 p0768 n0768 0 tlump
xseg0768 p0768 n0768 p0769 n0769 0 tlump
xseg0769 p0769 n0769 p0770 n0770 0 tlump
xseg0770 p0770 n0770 p0771 n0771 0 tlump
xseg0771 p0771 n0771 p0772 n0772 0 tlump
xseg0772 p0772 n0772 p0773 n0773 0 tlump
xseg0773 p0773 n0773 p0774 n0774 0 tlump
xseg0774 p0774 n0774 p0775 n0775 0 tlump
xseg0775 p0775 n0775 p0776 n0776 0 tlump
xseg0776 p0776 n0776 p0777 n0777 0 tlump
xseg0777 p0777 n0777 p0778 n0778 0 tlump
xseg0778 p0778 n0778 p0779 n0779 0 tlump
xseg0779 p0779 n0779 p0780 n0780 0 tlump
xseg0780 p0780 n0780 p0781 n0781 0 tlump
xseg0781 p0781 n0781 p0782 n0782 0 tlump
xseg0782 p0782 n0782 p0783 n0783 0 tlump
xseg0783 p0783 n0783 p0784 n0784 0 tlump
xseg0784 p0784 n0784 p0785 n0785 0 tlump
xseg0785 p0785 n0785 p0786 n0786 0 tlump
xseg0786 p0786 n0786 p0787 n0787 0 tlump
xseg0787 p0787 n0787 p0788 n0788 0 tlump
xseg0788 p0788 n0788 p0789 n0789 0 tlump
xseg0789 p0789 n0789 p0790 n0790 0 tlump
xseg0790 p0790 n0790 p0791 n0791 0 tlump
xseg0791 p0791 n0791 p0792 n0792 0 tlump
xseg0792 p0792 n0792 p0793 n0793 0 tlump
xseg0793 p0793 n0793 p0794 n0794 0 tlump
xseg0794 p0794 n0794 p0795 n0795 0 tlump
xseg0795 p0795 n0795 p0796 n0796 0 tlump
xseg0796 p0796 n0796 p0797 n0797 0 tlump
xseg0797 p0797 n0797 p0798 n0798 0 tlump
xseg0798 p0798 n0798 p0799 n0799 0 tlump
xseg0799 p0799 n0799 p0800 n0800 0 tlump
xseg0800 p0800 n0800 p0801 n0801 0 tlump
xseg0801 p0801 n0801 p0802 n0802 0 tlump
xseg0802 p0802 n0802 p0803 n0803 0 tlump
xseg0803 p0803 n0803 p0804 n0804 0 tlump
xseg0804 p0804 n0804 p0805 n0805 0 tlump
xseg0805 p0805 n0805 p0806 n0806 0 tlump
xseg0806 p0806 n0806 p0807 n0807 0 tlump
xseg0807 p0807 n0807 p0808 n0808 0 tlump
xseg0808 p0808 n0808 p0809 n0809 0 tlump
xseg0809 p0809 n0809 p0810 n0810 0 tlump
xseg0810 p0810 n0810 p0811 n0811 0 tlump
xseg0811 p0811 n0811 p0812 n0812 0 tlump
xseg0812 p0812 n0812 p0813 n0813 0 tlump
xseg0813 p0813 n0813 p0814 n0814 0 tlump
xseg0814 p0814 n0814 p0815 n0815 0 tlump
xseg0815 p0815 n0815 p0816 n0816 0 tlump
xseg0816 p0816 n0816 p0817 n0817 0 tlump
xseg0817 p0817 n0817 p0818 n0818 0 tlump
xseg0818 p0818 n0818 p0819 n0819 0 tlump
xseg0819 p0819 n0819 p0820 n0820 0 tlump
xseg0820 p0820 n0820 p0821 n0821 0 tlump
xseg0821 p0821 n0821 p0822 n0822 0 tlump
xseg0822 p0822 n0822 p0823 n0823 0 tlump
xseg0823 p0823 n0823 p0824 n0824 0 tlump
xseg0824 p0824 n0824 p0825 n0825 0 tlump
xseg0825 p0825 n0825 p0826 n0826 0 tlump
xseg0826 p0826 n0826 p0827 n0827 0 tlump
xseg0827 p0827 n0827 p0828 n0828 0 tlump
xseg0828 p0828 n0828 p0829 n0829 0 tlump
xseg0829 p0829 n0829 p0830 n0830 0 tlump
xseg0830 p0830 n0830 p0831 n0831 0 tlump
xseg0831 p0831 n0831 p0832 n0832 0 tlump
xseg0832 p0832 n0832 p0833 n0833 0 tlump
xseg0833 p0833 n0833 p0834 n0834 0 tlump
xseg0834 p0834 n0834 p0835 n0835 0 tlump
xseg0835 p0835 n0835 p0836 n0836 0 tlump
xseg0836 p0836 n0836 p0837 n0837 0 tlump
xseg0837 p0837 n0837 p0838 n0838 0 tlump
xseg0838 p0838 n0838 p0839 n0839 0 tlump
xseg0839 p0839 n0839 p0840 n0840 0 tlump
xseg0840 p0840 n0840 p0841 n0841 0 tlump
xseg0841 p0841 n0841 p0842 n0842 0 tlump
xseg0842 p0842 n0842 p0843 n0843 0 tlump
xseg0843 p0843 n0843 p0844 n0844 0 tlump
xseg0844 p0844 n0844 p0845 n0845 0 tlump
xseg0845 p0845 n0845 p0846 n0846 0 tlump
xseg0846 p0846 n0846 p0847 n0847 0 tlump
xseg0847 p0847 n0847 p0848 n0848 0 tlump
xseg0848 p0848 n0848 p0849 n0849 0 tlump
xseg0849 p0849 n0849 p0850 n0850 0 tlump
xseg0850 p0850 n0850 p0851 n0851 0 tlump
xseg0851 p0851 n0851 p0852 n0852 0 tlump
xseg0852 p0852 n0852 p0853 n0853 0 tlump
xseg0853 p0853 n0853 p0854 n0854 0 tlump
xseg0854 p0854 n0854 p0855 n0855 0 tlump
xseg0855 p0855 n0855 p0856 n0856 0 tlump
xseg0856 p0856 n0856 p0857 n0857 0 tlump
xseg0857 p0857 n0857 p0858 n0858 0 tlump
xseg0858 p0858 n0858 p0859 n0859 0 tlump
xseg0859 p0859 n0859 p0860 n0860 0 tlump
xseg0860 p0860 n0860 p0861 n0861 0 tlump
xseg0861 p0861 n0861 p0862 n0862 0 tlump
xseg0862 p0862 n0862 p0863 n0863 0 tlump
xseg0863 p0863 n0863 p0864 n0864 0 tlump
xseg0864 p0864 n0864 p0865 n0865 0 tlump
xseg0865 p0865 n0865 p0866 n0866 0 tlump
xseg0866 p0866 n0866 p0867 n0867 0 tlump
xseg0867 p0867 n0867 p0868 n0868 0 tlump
xseg0868 p0868 n0868 p0869 n0869 0 tlump
xseg0869 p0869 n0869 p0870 n0870 0 tlump
xseg0870 p0870 n0870 p0871 n0871 0 tlump
xseg0871 p0871 n0871 p0872 n0872 0 tlump
xseg0872 p0872 n0872 p0873 n0873 0 tlump
xseg0873 p0873 n0873 p0874 n0874 0 tlump
xseg0874 p0874 n0874 p0875 n0875 0 tlump
xseg0875 p0875 n0875 p0876 n0876 0 tlump
xseg0876 p0876 n0876 p0877 n0877 0 tlump
xseg0877 p0877 n0877 p0878 n0878 0 tlump
xseg0878 p0878 n0878 p0879 n0879 0 tlump
xseg0879 p0879 n0879 p0880 n0880 0 tlump
xseg0880 p0880 n0880 p0881 n0881 0 tlump
xseg0881 p0881 n0881 p0882 n0882 0 tlump
xseg0882 p0882 n0882 p0883 n0883 0 tlump
xseg0883 p0883 n0883 p0884 n0884 0 tlump
xseg0884 p0884 n0884 p0885 n0885 0 tlump
xseg0885 p0885 n0885 p0886 n0886 0 tlump
xseg0886 p0886 n0886 p0887 n0887 0 tlump
xseg0887 p0887 n0887 p0888 n0888 0 tlump
xseg0888 p0888 n0888 p0889 n0889 0 tlump
xseg0889 p0889 n0889 p0890 n0890 0 tlump
xseg0890 p0890 n0890 p0891 n0891 0 tlump
xseg0891 p0891 n0891 p0892 n0892 0 tlump
xseg0892 p0892 n0892 p0893 n0893 0 tlump
xseg0893 p0893 n0893 p0894 n0894 0 tlump
xseg0894 p0894 n0894 p0895 n0895 0 tlump
xseg0895 p0895 n0895 p0896 n0896 0 tlump
xseg0896 p0896 n0896 p0897 n0897 0 tlump
xseg0897 p0897 n0897 p0898 n0898 0 tlump
xseg0898 p0898 n0898 p0899 n0899 0 tlump
xseg0899 p0899 n0899 p0900 n0900 0 tlump
xseg0900 p0900 n0900 p0901 n0901 0 tlump
xseg0901 p0901 n0901 p0902 n0902 0 tlump
xseg0902 p0902 n0902 p0903 n0903 0 tlump
xseg0903 p0903 n0903 p0904 n0904 0 tlump
xseg0904 p0904 n0904 p0905 n0905 0 tlump
xseg0905 p0905 n0905 p0906 n0906 0 tlump
xseg0906 p0906 n0906 p0907 n0907 0 tlump
xseg0907 p0907 n0907 p0908 n0908 0 tlump
xseg0908 p0908 n0908 p0909 n0909 0 tlump
xseg0909 p0909 n0909 p0910 n0910 0 tlump
xseg0910 p0910 n0910 p0911 n0911 0 tlump
xseg0911 p0911 n0911 p0912 n0912 0 tlump
xseg0912 p0912 n0912 p0913 n0913 0 tlump
xseg0913 p0913 n0913 p0914 n0914 0 tlump
xseg0914 p0914 n0914 p0915 n0915 0 tlump
xseg0915 p0915 n0915 p0916 n0916 0 tlump
xseg0916 p0916 n0916 p0917 n0917 0 tlump
xseg0917 p0917 n0917 p0918 n0918 0 tlump
xseg0918 p0918 n0918 p0919 n0919 0 tlump
xseg0919 p0919 n0919 p0920 n0920 0 tlump
xseg0920 p0920 n0920 p0921 n0921 0 tlump
xseg0921 p0921 n0921 p0922 n0922 0 tlump
xseg0922 p0922 n0922 p0923 n0923 0 tlump
xseg0923 p0923 n0923 p0924 n0924 0 tlump
xseg0924 p0924 n0924 p0925 n0925 0 tlump
xseg0925 p0925 n0925 p0926 n0926 0 tlump
xseg0926 p0926 n0926 p0927 n0927 0 tlump
xseg0927 p0927 n0927 p0928 n0928 0 tlump
xseg0928 p0928 n0928 p0929 n0929 0 tlump
xseg0929 p0929 n0929 p0930 n0930 0 tlump
xseg0930 p0930 n0930 p0931 n0931 0 tlump
xseg0931 p0931 n0931 p0932 n0932 0 tlump
xseg0932 p0932 n0932 p0933 n0933 0 tlump
xseg0933 p0933 n0933 p0934 n0934 0 tlump
xseg0934 p0934 n0934 p0935 n0935 0 tlump
xseg0935 p0935 n0935 p0936 n0936 0 tlump
xseg0936 p0936 n0936 p0937 n0937 0 tlump
xseg0937 p0937 n0937 p0938 n0938 0 tlump
xseg0938 p0938 n0938 p0939 n0939 0 tlump
xseg0939 p0939 n0939 p0940 n0940 0 tlump
xseg0940 p0940 n0940 p0941 n0941 0 tlump
xseg0941 p0941 n0941 p0942 n0942 0 tlump
xseg0942 p0942 n0942 p0943 n0943 0 tlump
xseg0943 p0943 n0943 p0944 n0944 0 tlump
xseg0944 p0944 n0944 p0945 n0945 0 tlump
xseg0945 p0945 n0945 p0946 n0946 0 tlump
xseg0946 p0946 n0946 p0947 n0947 0 tlump
xseg0947 p0947 n0947 p0948 n0948 0 tlump
xseg0948 p0948 n0948 p0949 n0949 0 tlump
xseg0949 p0949 n0949 p0950 n0950 0 tlump
xseg0950 p0950 n0950 p0951 n0951 0 tlump
xseg0951 p0951 n0951 p0952 n0952 0 tlump
xseg0952 p0952 n0952 p0953 n0953 0 tlump
xseg0953 p0953 n0953 p0954 n0954 0 tlump
xseg0954 p0954 n0954 p0955 n0955 0 tlump
xseg0955 p0955 n0955 p0956 n0956 0 tlump
xseg0956 p0956 n0956 p0957 n0957 0 tlump
xseg0957 p0957 n0957 p0958 n0958 0 tlump
xseg0958 p0958 n0958 p0959 n0959 0 tlump
xseg0959 p0959 n0959 p0960 n0960 0 tlump
xseg0960 p0960 n0960 p0961 n0961 0 tlump
xseg0961 p0961 n0961 p0962 n0962 0 tlump
xseg0962 p0962 n0962 p0963 n0963 0 tlump
xseg0963 p0963 n0963 p0964 n0964 0 tlump
xseg0964 p0964 n0964 p0965 n0965 0 tlump
xseg0965 p0965 n0965 p0966 n0966 0 tlump
xseg0966 p0966 n0966 p0967 n0967 0 tlump
xseg0967 p0967 n0967 p0968 n0968 0 tlump
xseg0968 p0968 n0968 p0969 n0969 0 tlump
xseg0969 p0969 n0969 p0970 n0970 0 tlump
xseg0970 p0970 n0970 p0971 n0971 0 tlump
xseg0971 p0971 n0971 p0972 n0972 0 tlump
xseg0972 p0972 n0972 p0973 n0973 0 tlump
xseg0973 p0973 n0973 p0974 n0974 0 tlump
xseg0974 p0974 n0974 p0975 n0975 0 tlump
xseg0975 p0975 n0975 p0976 n0976 0 tlump
xseg0976 p0976 n0976 p0977 n0977 0 tlump
xseg0977 p0977 n0977 p0978 n0978 0 tlump
xseg0978 p0978 n0978 p0979 n0979 0 tlump
xseg0979 p0979 n0979 p0980 n0980 0 tlump
xseg0980 p0980 n0980 p0981 n0981 0 tlump
xseg0981 p0981 n0981 p0982 n0982 0 tlump
xseg0982 p0982 n0982 p0983 n0983 0 tlump
xseg0983 p0983 n0983 p0984 n0984 0 tlump
xseg0984 p0984 n0984 p0985 n0985 0 tlump
xseg0985 p0985 n0985 p0986 n0986 0 tlump
xseg0986 p0986 n0986 p0987 n0987 0 tlump
xseg0987 p0987 n0987 p0988 n0988 0 tlump
xseg0988 p0988 n0988 p0989 n0989 0 tlump
xseg0989 p0989 n0989 p0990 n0990 0 tlump
xseg0990 p0990 n0990 p0991 n0991 0 tlump
xseg0991 p0991 n0991 p0992 n0992 0 tlump
xseg0992 p0992 n0992 p0993 n0993 0 tlump
xseg0993 p0993 n0993 p0994 n0994 0 tlump
xseg0994 p0994 n0994 p0995 n0995 0 tlump
xseg0995 p0995 n0995 p0996 n0996 0 tlump
xseg0996 p0996 n0996 p0997 n0997 0 tlump
xseg0997 p0997 n0997 p0998 n0998 0 tlump
xseg0998 p0998 n0998 p0999 n0999 0 tlump
xseg0999 p0999 n0999 p1000 n1000 0 tlump
rend_term p1000 n1000 100.000000
**************************
***** pd attachments *****
**************************
*pd 01 - attach at 0.000 meters with 0.000 meter drop
xseg0012_0000 p0012 n0012 p0012_0001 n0012_0001 0 tlump
xseg0012_0001 p0012_0001 n0012_0001 p0012_0002 n0012_0002 0 tlump
xseg0012_0002 p0012_0002 n0012_0002 p0012_0003 n0012_0003 0 tlump
xseg0012_0003 p0012_0003 n0012_0003 p0012_0004 n0012_0004 0 tlump
xseg0012_0004 p0012_0004 n0012_0004 p0012_0005 n0012_0005 0 tlump
xseg0012_0005 p0012_0005 n0012_0005 p0012_0006 n0012_0006 0 tlump
rpdp0012 p0012_0006 pdp_0001 0.010
rpdn0012 n0012_0006 pdn_0001 0.010
xpd0001 pdp_0001 pdn_0001 0 pd
*pd 02 - attach at 41.000 meters with 0.000 meter drop
xseg0832_0000 p0832 n0832 p0832_0001 n0832_0001 0 tlump
xseg0832_0001 p0832_0001 n0832_0001 p0832_0002 n0832_0002 0 tlump
xseg0832_0002 p0832_0002 n0832_0002 p0832_0003 n0832_0003 0 tlump
xseg0832_0003 p0832_0003 n0832_0003 p0832_0004 n0832_0004 0 tlump
xseg0832_0004 p0832_0004 n0832_0004 p0832_0005 n0832_0005 0 tlump
xseg0832_0005 p0832_0005 n0832_0005 p0832_0006 n0832_0006 0 tlump
rpdp0832 p0832_0006 pdp_0002 0.010
rpdn0832 n0832_0006 pdn_0002 0.010
xpd0002 pdp_0002 pdn_0002 0 pd
*pd 03 - attach at 42.000 meters with 0.000 meter drop
xseg0844_0000 p0844 n0844 p0844_0001 n0844_0001 0 tlump
xseg0844_0001 p0844_0001 n0844_0001 p0844_0002 n0844_0002 0 tlump
xseg0844_0002 p0844_0002 n0844_0002 p0844_0003 n0844_0003 0 tlump
xseg0844_0003 p0844_0003 n0844_0003 p0844_0004 n0844_0004 0 tlump
xseg0844_0004 p0844_0004 n0844_0004 p0844_0005 n0844_0005 0 tlump
xseg0844_0005 p0844_0005 n0844_0005 p0844_0006 n0844_0006 0 tlump
rpdp0844 p0844_0006 pdp_0003 0.010
rpdn0844 n0844_0006 pdn_0003 0.010
xpd0003 pdp_0003 pdn_0003 0 pd
vac p0000_p n0000_n 0 ac 1
rp p0000 p0000_p 50
rn n0000_n n0000 50
rrpp p0000_p refp 50
rrpn refp 0 50
rrnp n0000_n refn 50
rrnn refn 0 50
.ac lin 500 1meg 100meg
.net i(rend_term) vac
.save  v(refp) v(refn)  i(vac) i(rp) i(rend_term)  v(p0000) v(n0000)  s11(vac) s21(vac)  v(p1000) v(n1000)
