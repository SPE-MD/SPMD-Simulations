*tranient sim command for cable impedance measurement
.include cable.p
vap ap 0 0
+pwl 0 0
++50n  0.0
++10n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++10n  0.0
van 0 an 0
+pwl 0 0
++50n  0.0
++10n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n -1.0
++20n  1.0
++20n  1.0
++10n  0.0
rap ap p0000 50
ran an n0000 50
rrefp ap refp 50
rrefn an refn 50
rref  refp refn 100
.save V(*)
.tran 2000n
